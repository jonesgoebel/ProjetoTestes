LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.numeric_std.all;


entity FMELUMA is
	port (
		CLK: IN std_logic;
		RESET: IN std_logic;		
		A0, A1, A2, A3, A4, A5, A6, A7, A8, A9, A10, A11, A12, A13, A14: IN std_logic_vector(7 downto 0);--AMOSTRAS PARA SEREM INTERPOLADAS
		B0, B1, B2, B3, B4, B5, B6, B7: IN std_logic_vector(7 downto 0);--AMOSTRAS ORIGINAIS PARA COMPARAÇÃO
		LOAD_A: OUT  std_logic;
		LOAD_B: OUT  std_logic;
		READY: OUT  std_logic;	
		MVX,MVY: OUT bit_vector(2 downto 0);
		SAD: OUT std_logic_vector(16 downto 0)
	);
end FMELUMA;

architecture arc of FMELUMA is
	
	SIGNAL S0,S1,S2,S3,S4,S5,S6,S7: std_logic_vector(11 downto 0);
	SIGNAL S8,S9,S10,S11,S12,S13,S14,S15: std_logic_vector(11 downto 0);
	SIGNAL S16,S17,S18,S19,S20,S21,S22,S23: std_logic_vector(11 downto 0);
	SIGNAL S24,S25,S26,S27,S28,S29,S30,S31: std_logic_vector(11 downto 0);
	SIGNAL S32,S33,S34,S35,S36,S37,S38,S39: std_logic_vector(11 downto 0);
	SIGNAL S40,S41,S42,S43,S44,S45,S46,S47: std_logic_vector(11 downto 0);
	SIGNAL S48,S49,S50,S51,S52,S53,S54,S55: std_logic_vector(11 downto 0);
	SIGNAL S56,S57,S58,S59,S60,S61,S62,S63: std_logic_vector(11 downto 0);
	SIGNAL S64,S65,S66,S67,S68,S69,S70,S71: std_logic_vector(11 downto 0);
	SIGNAL S72,S73,S74,S75,S76,S77,S78,S79: std_logic_vector(11 downto 0);
	SIGNAL S80,S81,S82,S83,S84,S85,S86,S87: std_logic_vector(11 downto 0);
	SIGNAL S88,S89,S90,S91,S92,S93,S94,S95: std_logic_vector(11 downto 0);
	SIGNAL S96,S97,S98,S99,S100,S101,S102,S103: std_logic_vector(11 downto 0);
	SIGNAL S104,S105,S106,S107,S108,S109,S110,S111: std_logic_vector(11 downto 0);
	SIGNAL S112,S113,S114,S115,S116,S117,S118,S119: std_logic_vector(11 downto 0);
	SIGNAL S120,S121,S122,S123,S124,S125,S126,S127: std_logic_vector(11 downto 0);
    SIGNAL S128,S129,S130,S131,S132,S133,S134,S135: std_logic_vector(11 downto 0);
    SIGNAL S136,S137,S138,S139,S140,S141,S142,S143: std_logic_vector(11 downto 0);
    SIGNAL S144,S145,S146,S147,S148,S149,S150,S151: std_logic_vector(11 downto 0);
    SIGNAL S152,S153,S154,S155,S156,S157,S158,S159: std_logic_vector(11 downto 0);
    SIGNAL S160,S161,S162,S163,S164,S165,S166,S167: std_logic_vector(11 downto 0);
    SIGNAL S168,S169,S170,S171,S172,S173,S174,S175: std_logic_vector(11 downto 0);
    SIGNAL S176,S177,S178,S179,S180,S181,S182,S183: std_logic_vector(11 downto 0);
    SIGNAL S184,S185,S186,S187,S188,S189,S190,S191: std_logic_vector(11 downto 0);
    SIGNAL S192,S193,S194,S195,S196,S197,S198,S199: std_logic_vector(11 downto 0);
    SIGNAL S200,S201,S202,S203,S204,S205,S206,S207: std_logic_vector(11 downto 0);
    SIGNAL S208,S209,S210,S211,S212,S213,S214,S215: std_logic_vector(11 downto 0);
    SIGNAL S216,S217,S218,S219,S220,S221,S222,S223: std_logic_vector(11 downto 0);
    SIGNAL S224,S225,S226,S227,S228,S229,S230,S231: std_logic_vector(11 downto 0);
    SIGNAL S232,S233,S234,S235,S236,S237,S238,S239: std_logic_vector(11 downto 0);
    SIGNAL S240,S241,S242,S243,S244,S245,S246,S247: std_logic_vector(11 downto 0);
    SIGNAL S248,S249,S250,S251,S252,S253,S254,S255: std_logic_vector(11 downto 0);
    SIGNAL S256,S257,S258,S259,S260,S261,S262,S263: std_logic_vector(11 downto 0);
    SIGNAL S264,S265,S266,S267,S268,S269,S270,S271: std_logic_vector(11 downto 0);
    SIGNAL S272,S273,S274,S275,S276,S277,S278,S279: std_logic_vector(11 downto 0);
    SIGNAL S280,S281,S282,S283,S284,S285,S286,S287: std_logic_vector(11 downto 0);
    SIGNAL S288,S289,S290,S291,S292,S293,S294,S295: std_logic_vector(11 downto 0);
    SIGNAL S296,S297,S298,S299,S300,S301,S302,S303: std_logic_vector(11 downto 0);
    SIGNAL S304,S305,S306,S307,S308,S309,S310,S311: std_logic_vector(11 downto 0);
    SIGNAL S312,S313,S314,S315,S316,S317,S318,S319: std_logic_vector(11 downto 0);
    SIGNAL S320,S321,S322,S323,S324,S325,S326,S327: std_logic_vector(11 downto 0);
    SIGNAL S328,S329,S330,S331,S332,S333,S334,S335: std_logic_vector(11 downto 0);
    SIGNAL S336,S337,S338,S339,S340,S341,S342,S343: std_logic_vector(11 downto 0);
    SIGNAL S344,S345,S346,S347,S348,S349,S350,S351: std_logic_vector(11 downto 0);
    SIGNAL S352,S353,S354,S355,S356,S357,S358,S359: std_logic_vector(11 downto 0);
    SIGNAL S360,S361,S362,S363,S364,S365,S366,S367: std_logic_vector(11 downto 0);
    SIGNAL S368,S369,S370,S371,S372,S373,S374,S375: std_logic_vector(11 downto 0);
    SIGNAL S376,S377,S378,S379,S380,S381,S382,S383: std_logic_vector(11 downto 0);
    SIGNAL S384,S385,S386,S387,S388,S389,S390,S391: std_logic_vector(11 downto 0);
    SIGNAL S392,S393,S394,S395,S396,S397,S398,S399: std_logic_vector(11 downto 0);
    SIGNAL S400,S401,S402,S403,S404,S405,S406,S407: std_logic_vector(11 downto 0);
    SIGNAL S408,S409,S410,S411,S412,S413,S414,S415: std_logic_vector(11 downto 0);
    SIGNAL S416,S417,S418,S419,S420,S421,S422,S423: std_logic_vector(11 downto 0);
    SIGNAL S424,S425,S426,S427,S428,S429,S430,S431: std_logic_vector(11 downto 0);
    SIGNAL S432,S433,S434,S435,S436,S437,S438,S439: std_logic_vector(11 downto 0);
    SIGNAL S440,S441,S442,S443,S444,S445,S446,S447: std_logic_vector(11 downto 0);
    SIGNAL S448,S449,S450,S451,S452,S453,S454,S455: std_logic_vector(11 downto 0);
    SIGNAL S456,S457,S458,S459,S460,S461,S462,S463: std_logic_vector(11 downto 0);
    SIGNAL S464,S465,S466,S467,S468,S469,S470,S471: std_logic_vector(11 downto 0);
    SIGNAL S472,S473,S474,S475,S476,S477,S478,S479: std_logic_vector(11 downto 0);
    SIGNAL S480,S481,S482,S483,S484,S485,S486,S487: std_logic_vector(11 downto 0);
    SIGNAL S488,S489,S490,S491,S492,S493,S494,S495: std_logic_vector(11 downto 0);
    SIGNAL S496,S497,S498,S499,S500,S501,S502,S503: std_logic_vector(11 downto 0);
    SIGNAL S504,S505,S506,S507,S508,S509,S510,S511: std_logic_vector(11 downto 0);
	
	
	
	SIGNAL 	R0,R1,R2,R3,R4,R5,R6,R7,R8,R9,R10,R11,R12,R13,R14,R15,
			R16,R17,R18,R19,R20,R21,R22,R23,R24,R25,R26,R27,R28,R29,R30,R31,
			R32,R33,R34,R35,R36,R37,R38,R39,R40,R41,R42,R43,R44,R45,R46,R47,
			R48,R49,R50,R51,R52,R53,R54,R55,R56,R57,R58,R59,R60,R61,R62,R63: std_logic_vector(11 downto 0);
	
	SIGNAL ENABLE_RI, RESET_SAD,ENABLE_SAD,RESET_BEST_SAD :std_logic;
	SIGNAL SELETOR :BIT_VECTOR(2 downto 0);
	
	COMPONENT LumaInterpolation IS
		port (
		CLK: IN std_logic;
		ENABLE: IN std_logic;		
		A0, A1, A2, A3, A4, A5, A6, A7, A8, A9, A10, A11, A12, A13, A14: IN std_logic_vector(7 downto 0);
		S0,S1,S2,S3,S4,S5,S6,S7: OUT std_logic_vector(11 downto 0);
		S8,S9,S10,S11,S12,S13,S14,S15: OUT std_logic_vector(11 downto 0);
		S16,S17,S18,S19,S20,S21,S22,S23: OUT std_logic_vector(11 downto 0);
		S24,S25,S26,S27,S28,S29,S30,S31: OUT std_logic_vector(11 downto 0);
		S32,S33,S34,S35,S36,S37,S38,S39: OUT std_logic_vector(11 downto 0);
		S40,S41,S42,S43,S44,S45,S46,S47: OUT std_logic_vector(11 downto 0);
		S48,S49,S50,S51,S52,S53,S54,S55: OUT std_logic_vector(11 downto 0);
		S56,S57,S58,S59,S60,S61,S62,S63: OUT std_logic_vector(11 downto 0);
		S64,S65,S66,S67,S68,S69,S70,S71: OUT std_logic_vector(11 downto 0);
		S72,S73,S74,S75,S76,S77,S78,S79: OUT std_logic_vector(11 downto 0);
		S80,S81,S82,S83,S84,S85,S86,S87: OUT std_logic_vector(11 downto 0);
		S88,S89,S90,S91,S92,S93,S94,S95: OUT std_logic_vector(11 downto 0);
		S96,S97,S98,S99,S100,S101,S102,S103: OUT std_logic_vector(11 downto 0);
		S104,S105,S106,S107,S108,S109,S110,S111: OUT std_logic_vector(11 downto 0);
		S112,S113,S114,S115,S116,S117,S118,S119: OUT std_logic_vector(11 downto 0);
		S120,S121,S122,S123,S124,S125,S126,S127: OUT std_logic_vector(11 downto 0);
        S128,S129,S130,S131,S132,S133,S134,S135: OUT std_logic_vector(11 downto 0);
        S136,S137,S138,S139,S140,S141,S142,S143: OUT std_logic_vector(11 downto 0);
        S144,S145,S146,S147,S148,S149,S150,S151: OUT std_logic_vector(11 downto 0);
        S152,S153,S154,S155,S156,S157,S158,S159: OUT std_logic_vector(11 downto 0);
        S160,S161,S162,S163,S164,S165,S166,S167: OUT std_logic_vector(11 downto 0);
        S168,S169,S170,S171,S172,S173,S174,S175: OUT std_logic_vector(11 downto 0);
        S176,S177,S178,S179,S180,S181,S182,S183: OUT std_logic_vector(11 downto 0);
        S184,S185,S186,S187,S188,S189,S190,S191: OUT std_logic_vector(11 downto 0);
        S192,S193,S194,S195,S196,S197,S198,S199: OUT std_logic_vector(11 downto 0);
        S200,S201,S202,S203,S204,S205,S206,S207: OUT std_logic_vector(11 downto 0);
        S208,S209,S210,S211,S212,S213,S214,S215: OUT std_logic_vector(11 downto 0);
        S216,S217,S218,S219,S220,S221,S222,S223: OUT std_logic_vector(11 downto 0);
        S224,S225,S226,S227,S228,S229,S230,S231: OUT std_logic_vector(11 downto 0);
        S232,S233,S234,S235,S236,S237,S238,S239: OUT std_logic_vector(11 downto 0);
        S240,S241,S242,S243,S244,S245,S246,S247: OUT std_logic_vector(11 downto 0);
        S248,S249,S250,S251,S252,S253,S254,S255: OUT std_logic_vector(11 downto 0);
        S256,S257,S258,S259,S260,S261,S262,S263: OUT std_logic_vector(11 downto 0);
        S264,S265,S266,S267,S268,S269,S270,S271: OUT std_logic_vector(11 downto 0);
        S272,S273,S274,S275,S276,S277,S278,S279: OUT std_logic_vector(11 downto 0);
        S280,S281,S282,S283,S284,S285,S286,S287: OUT std_logic_vector(11 downto 0);
        S288,S289,S290,S291,S292,S293,S294,S295: OUT std_logic_vector(11 downto 0);
        S296,S297,S298,S299,S300,S301,S302,S303: OUT std_logic_vector(11 downto 0);
        S304,S305,S306,S307,S308,S309,S310,S311: OUT std_logic_vector(11 downto 0);
        S312,S313,S314,S315,S316,S317,S318,S319: OUT std_logic_vector(11 downto 0);
        S320,S321,S322,S323,S324,S325,S326,S327: OUT std_logic_vector(11 downto 0);
        S328,S329,S330,S331,S332,S333,S334,S335: OUT std_logic_vector(11 downto 0);
        S336,S337,S338,S339,S340,S341,S342,S343: OUT std_logic_vector(11 downto 0);
        S344,S345,S346,S347,S348,S349,S350,S351: OUT std_logic_vector(11 downto 0);
        S352,S353,S354,S355,S356,S357,S358,S359: OUT std_logic_vector(11 downto 0);
        S360,S361,S362,S363,S364,S365,S366,S367: OUT std_logic_vector(11 downto 0);
        S368,S369,S370,S371,S372,S373,S374,S375: OUT std_logic_vector(11 downto 0);
        S376,S377,S378,S379,S380,S381,S382,S383: OUT std_logic_vector(11 downto 0);
        S384,S385,S386,S387,S388,S389,S390,S391: OUT std_logic_vector(11 downto 0);
        S392,S393,S394,S395,S396,S397,S398,S399: OUT std_logic_vector(11 downto 0);
        S400,S401,S402,S403,S404,S405,S406,S407: OUT std_logic_vector(11 downto 0);
        S408,S409,S410,S411,S412,S413,S414,S415: OUT std_logic_vector(11 downto 0);
        S416,S417,S418,S419,S420,S421,S422,S423: OUT std_logic_vector(11 downto 0);
        S424,S425,S426,S427,S428,S429,S430,S431: OUT std_logic_vector(11 downto 0);
        S432,S433,S434,S435,S436,S437,S438,S439: OUT std_logic_vector(11 downto 0);
        S440,S441,S442,S443,S444,S445,S446,S447: OUT std_logic_vector(11 downto 0);
        S448,S449,S450,S451,S452,S453,S454,S455: OUT std_logic_vector(11 downto 0);
        S456,S457,S458,S459,S460,S461,S462,S463: OUT std_logic_vector(11 downto 0);
        S464,S465,S466,S467,S468,S469,S470,S471: OUT std_logic_vector(11 downto 0);
        S472,S473,S474,S475,S476,S477,S478,S479: OUT std_logic_vector(11 downto 0);
        S480,S481,S482,S483,S484,S485,S486,S487: OUT std_logic_vector(11 downto 0);
        S488,S489,S490,S491,S492,S493,S494,S495: OUT std_logic_vector(11 downto 0);
        S496,S497,S498,S499,S500,S501,S502,S503: OUT std_logic_vector(11 downto 0);
        S504,S505,S506,S507,S508,S509,S510,S511: OUT std_logic_vector(11 downto 0)
	);
	END COMPONENT;	
		
	COMPONENT Arvore_sad IS
		port (
			S0,S1,S2,S3,S4,S5,S6,S7: IN std_logic_vector(11 downto 0);
			S8,S9,S10,S11,S12,S13,S14,S15: IN std_logic_vector(11 downto 0);
			S16,S17,S18,S19,S20,S21,S22,S23: IN std_logic_vector(11 downto 0);
			S24,S25,S26,S27,S28,S29,S30,S31: IN std_logic_vector(11 downto 0);
			S32,S33,S34,S35,S36,S37,S38,S39: IN std_logic_vector(11 downto 0);
			S40,S41,S42,S43,S44,S45,S46,S47: IN std_logic_vector(11 downto 0);
			S48,S49,S50,S51,S52,S53,S54,S55: IN std_logic_vector(11 downto 0);
			S56,S57,S58,S59,S60,S61,S62,S63: IN std_logic_vector(11 downto 0);
			b0,b1,b2,b3,b4,b5,b6,b7 : in  std_logic_vector(7 downto 0);
			r0,r1,r2,r3,r4,r5,r6,r7 : out std_logic_vector(11 downto 0)
		);
	END COMPONENT;
	
	COMPONENT SAD_reg is
		port (
			CLK: IN std_logic;
			RESET_SAD: IN std_logic;
			ENABLE_SAD: IN std_logic;
			SELETOR: IN BIT_VECTOR(2 downto 0);
			RESET_BEST_SAD: IN std_logic;	
			A0,A1,A2,A3,A4,A5,A6,A7,A8,A9,A10,A11,A12,A13,A14,A15,
			A16,A17,A18,A19,A20,A21,A22,A23,A24,A25,A26,A27,A28,A29,A30,A31,
			A32,A33,A34,A35,A36,A37,A38,A39,A40,A41,A42,A43,A44,A45,A46,A47,
			A48,A49,A50,A51,A52,A53,A54,A55,A56,A57,A58,A59,A60,A61,A62,A63: IN std_logic_vector(11 downto 0);
			MVX,MVY: OUT bit_vector(2 downto 0);
			SAD: OUT std_logic_vector(16 downto 0)
		);
	END COMPONENT;
	
	COMPONENT controle is
		port (
			CLK: IN std_logic;
			RESET: IN std_logic;
			READY: OUT  std_logic;	
			LOAD_A: OUT  std_logic;
			LOAD_B: OUT  std_logic;
			ENABLE_RI: OUT  std_logic;	
			SELETOR: OUT BIT_VECTOR(2 downto 0);
			RESET_SAD: OUT std_logic;
			ENABLE_SAD: OUT std_logic;
			RESET_BEST_SAD: OUT std_logic
		);
	END COMPONENT;
	
begin
	Inter: LumaInterpolation port map(CLK,ENABLE_RI,A0, A1, A2, A3, A4, A5, A6, A7, A8, A9, A10, A11, A12, A13, A14,
					S0,S1,S2,S3,S4,S5,S6,S7,S8,S9,S10,S11,S12,S13,S14,S15,
					S16,S17,S18,S19,S20,S21,S22,S23,S24,S25,S26,S27,S28,S29,S30,S31,
					S32,S33,S34,S35,S36,S37,S38,S39,S40,S41,S42,S43,S44,S45,S46,S47,
					S48,S49,S50,S51,S52,S53,S54,S55,S56,S57,S58,S59,S60,S61,S62,S63,
					S64,S65,S66,S67,S68,S69,S70,S71,S72,S73,S74,S75,S76,S77,S78,S79,
					S80,S81,S82,S83,S84,S85,S86,S87,S88,S89,S90,S91,S92,S93,S94,S95,
					S96,S97,S98,S99,S100,S101,S102,S103,S104,S105,S106,S107,S108,S109,S110,S111,
					S112,S113,S114,S115,S116,S117,S118,S119,S120,S121,S122,S123,S124,S125,S126,S127,
					S128,S129,S130,S131,S132,S133,S134,S135,S136,S137,S138,S139,S140,S141,S142,S143,
					S144,S145,S146,S147,S148,S149,S150,S151,S152,S153,S154,S155,S156,S157,S158,S159,
					S160,S161,S162,S163,S164,S165,S166,S167,S168,S169,S170,S171,S172,S173,S174,S175,
					S176,S177,S178,S179,S180,S181,S182,S183,S184,S185,S186,S187,S188,S189,S190,S191,
					S192,S193,S194,S195,S196,S197,S198,S199,S200,S201,S202,S203,S204,S205,S206,S207,
					S208,S209,S210,S211,S212,S213,S214,S215,S216,S217,S218,S219,S220,S221,S222,S223,
					S224,S225,S226,S227,S228,S229,S230,S231,S232,S233,S234,S235,S236,S237,S238,S239,
					S240,S241,S242,S243,S244,S245,S246,S247,S248,S249,S250,S251,S252,S253,S254,S255,
					S256,S257,S258,S259,S260,S261,S262,S263,S264,S265,S266,S267,S268,S269,S270,S271,
					S272,S273,S274,S275,S276,S277,S278,S279,S280,S281,S282,S283,S284,S285,S286,S287,
					S288,S289,S290,S291,S292,S293,S294,S295,S296,S297,S298,S299,S300,S301,S302,S303,
					S304,S305,S306,S307,S308,S309,S310,S311,S312,S313,S314,S315,S316,S317,S318,S319,
					S320,S321,S322,S323,S324,S325,S326,S327,S328,S329,S330,S331,S332,S333,S334,S335,
					S336,S337,S338,S339,S340,S341,S342,S343,S344,S345,S346,S347,S348,S349,S350,S351,
					S352,S353,S354,S355,S356,S357,S358,S359,S360,S361,S362,S363,S364,S365,S366,S367,
					S368,S369,S370,S371,S372,S373,S374,S375,S376,S377,S378,S379,S380,S381,S382,S383,
					S384,S385,S386,S387,S388,S389,S390,S391,S392,S393,S394,S395,S396,S397,S398,S399,
					S400,S401,S402,S403,S404,S405,S406,S407,S408,S409,S410,S411,S412,S413,S414,S415,
					S416,S417,S418,S419,S420,S421,S422,S423,S424,S425,S426,S427,S428,S429,S430,S431,
					S432,S433,S434,S435,S436,S437,S438,S439,S440,S441,S442,S443,S444,S445,S446,S447,
					S448,S449,S450,S451,S452,S453,S454,S455,S456,S457,S458,S459,S460,S461,S462,S463,
					S464,S465,S466,S467,S468,S469,S470,S471,S472,S473,S474,S475,S476,S477,S478,S479,
					S480,S481,S482,S483,S484,S485,S486,S487,S488,S489,S490,S491,S492,S493,S494,S495,
					S496,S497,S498,S499,S500,S501,S502,S503,S504,S505,S506,S507,S508,S509,S510,S511);
					
	arvore_0: arvore_sad port map(S0,S1,S2,S3,S4,S5,S6,S7,S8,S9,S10,S11,S12,S13,S14,S15,
					S16,S17,S18,S19,S20,S21,S22,S23,S24,S25,S26,S27,S28,S29,S30,S31,
					S32,S33,S34,S35,S36,S37,S38,S39,S40,S41,S42,S43,S44,S45,S46,S47,
					S48,S49,S50,S51,S52,S53,S54,S55,S56,S57,S58,S59,S60,S61,S62,S63,
					B0,B1,B2,B3,B4,B5,B6,B7, R0,R1,R2,R3,R4,R5,R6,R7);
					
					
	arvore_1: arvore_sad port map(
					S64,S65,S66,S67,S68,S69,S70,S71,S72,S73,S74,S75,S76,S77,S78,S79,
					S80,S81,S82,S83,S84,S85,S86,S87,S88,S89,S90,S91,S92,S93,S94,S95,
					S96,S97,S98,S99,S100,S101,S102,S103,S104,S105,S106,S107,S108,S109,S110,S111,
					S112,S113,S114,S115,S116,S117,S118,S119,S120,S121,S122,S123,S124,S125,S126,S127,
					B0,B1,B2,B3,B4,B5,B6,B7, R8,R9,R10,R11,R12,R13,R14,R15);				
	
	arvore_2: arvore_sad port map(
					S128,S129,S130,S131,S132,S133,S134,S135,S136,S137,S138,S139,S140,S141,S142,S143,
					S144,S145,S146,S147,S148,S149,S150,S151,S152,S153,S154,S155,S156,S157,S158,S159,
					S160,S161,S162,S163,S164,S165,S166,S167,S168,S169,S170,S171,S172,S173,S174,S175,
					S176,S177,S178,S179,S180,S181,S182,S183,S184,S185,S186,S187,S188,S189,S190,S191,
					B0,B1,B2,B3,B4,B5,B6,B7, R16,R17,R18,R19,R20,R21,R22,R23);				
	
	arvore_3: arvore_sad port map(
					S192,S193,S194,S195,S196,S197,S198,S199,S200,S201,S202,S203,S204,S205,S206,S207,
					S208,S209,S210,S211,S212,S213,S214,S215,S216,S217,S218,S219,S220,S221,S222,S223,
					S224,S225,S226,S227,S228,S229,S230,S231,S232,S233,S234,S235,S236,S237,S238,S239,
					S240,S241,S242,S243,S244,S245,S246,S247,S248,S249,S250,S251,S252,S253,S254,S255,
					B0,B1,B2,B3,B4,B5,B6,B7, R24,R25,R26,R27,R28,R29,R30,R31);				
	
	arvore_4: arvore_sad port map(
					S256,S257,S258,S259,S260,S261,S262,S263,S264,S265,S266,S267,S268,S269,S270,S271,
					S272,S273,S274,S275,S276,S277,S278,S279,S280,S281,S282,S283,S284,S285,S286,S287,
					S288,S289,S290,S291,S292,S293,S294,S295,S296,S297,S298,S299,S300,S301,S302,S303,
					S304,S305,S306,S307,S308,S309,S310,S311,S312,S313,S314,S315,S316,S317,S318,S319,
					B0,B1,B2,B3,B4,B5,B6,B7, R32,R33,R34,R35,R36,R37,R38,R39);				
	
	arvore_5: arvore_sad port map(
					S320,S321,S322,S323,S324,S325,S326,S327,S328,S329,S330,S331,S332,S333,S334,S335,
					S336,S337,S338,S339,S340,S341,S342,S343,S344,S345,S346,S347,S348,S349,S350,S351,
					S352,S353,S354,S355,S356,S357,S358,S359,S360,S361,S362,S363,S364,S365,S366,S367,
					S368,S369,S370,S371,S372,S373,S374,S375,S376,S377,S378,S379,S380,S381,S382,S383,
					B0,B1,B2,B3,B4,B5,B6,B7, R40,R41,R42,R43,R44,R45,R46,R47);				
	
	arvore_6: arvore_sad port map(
					S384,S385,S386,S387,S388,S389,S390,S391,S392,S393,S394,S395,S396,S397,S398,S399,
					S400,S401,S402,S403,S404,S405,S406,S407,S408,S409,S410,S411,S412,S413,S414,S415,
					S416,S417,S418,S419,S420,S421,S422,S423,S424,S425,S426,S427,S428,S429,S430,S431,
					S432,S433,S434,S435,S436,S437,S438,S439,S440,S441,S442,S443,S444,S445,S446,S447,
					B0,B1,B2,B3,B4,B5,B6,B7, R48,R49,R50,R51,R52,R53,R54,R55);				
	
	arvore_7: arvore_sad port map(
					S448,S449,S450,S451,S452,S453,S454,S455,S456,S457,S458,S459,S460,S461,S462,S463,
					S464,S465,S466,S467,S468,S469,S470,S471,S472,S473,S474,S475,S476,S477,S478,S479,
					S480,S481,S482,S483,S484,S485,S486,S487,S488,S489,S490,S491,S492,S493,S494,S495,
					S496,S497,S498,S499,S500,S501,S502,S503,S504,S505,S506,S507,S508,S509,S510,S511,
					B0,B1,B2,B3,B4,B5,B6,B7, R56,R57,R58,R59,R60,R61,R62,R63);				
	
	
	result_sad: SAD_reg port map(CLK,RESET_SAD,ENABLE_SAD,SELETOR,RESET_BEST_SAD,
								R0,R1,R2,R3,R4,R5,R6,R7,R8,R9,R10,R11,R12,R13,R14,R15,
								R16,R17,R18,R19,R20,R21,R22,R23,R24,R25,R26,R27,R28,R29,R30,R31,
								R32,R33,R34,R35,R36,R37,R38,R39,R40,R41,R42,R43,R44,R45,R46,R47,
								R48,R49,R50,R51,R52,R53,R54,R55,R56,R57,R58,R59,R60,R61,R62,R63,
								MVY,MVX,SAD);
					
	control: controle port map(CLK,RESET,READY,LOAD_A,LOAD_B,ENABLE_RI,SELETOR,
									RESET_SAD,ENABLE_SAD,RESET_BEST_SAD);
				
	
end arc;
